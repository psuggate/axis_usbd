`timescale 1ns / 100ps
module axis_usbd_tb;

endmodule // axis_usbd_tb
